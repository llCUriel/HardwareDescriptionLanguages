LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Hw3 IS

	PORT(
		 A : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		 B : IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Ax: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 By: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 test: OUT STD_LOGIC
		);

END Hw3;

ARCHITECTURE Hw3Architecture OF Hw3 IS

BEGIN
	PROCESS(A,B,Test)
	BEGIN
		IF(Test ='1') THEN
			Ax<= A and B;
		ELSIF(Test = '0') THEN
			By<= A or B;
		END IF;
	END PROCESS;
END Hw3Architecture;
