LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_BIT.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY Mux IS
	PORT (
		A	  : IN  STD_LOGIC;
		B    : IN  STD_LOGIC;
		C	  : OUT STD_LOGIC;
		S    : IN STD_LOGIC
	);
 
END Mux;

ARCHITECTURE MuxA OF Mux IS

BEGIN

	C <= A when S else B;
	
END MuxA;