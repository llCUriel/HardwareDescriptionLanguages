LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_BIT.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY Multiplexer_2_To_1T IS
	PORT (
		A	  : IN  STD_LOGIC_VECTOR(6 DOWNTO 0);
		B    : IN  STD_LOGIC_VECTOR(6 DOWNTO 0);
		C	  : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		S    : IN STD_LOGIC
	);
 
END Multiplexer_2_To_1T;

ARCHITECTURE MuxA OF Multiplexer_2_To_1T IS

BEGIN

	C <= B when S else A;
	
END MuxA;