LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Hw3 IS

	PORT(
		 DATA_IN : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		 SHAMNT  : IN 	STD_LOGIC_VECTOR(2 DOWNTO 0);
		 DATA_OUT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);

END Hw3;

ARCHITECTURE Hw3Architecture OF Hw3 IS

BEGIN
	PROCESS(DATA_IN,SHAMNT)
	BEGIN
		CASE SHAMNT IS
			WHEN "001"  => DATA_OUT <= '0' & DATA_IN(3 DOWNTO 1);
			WHEN "010"  => DATA_OUT <= DATA_IN(2 DOWNTO 0) & '0';
			WHEN "011"  => DATA_OUT <= DATA_IN(0) & DATA_IN(3 DOWNTO 1);
			WHEN "100"  => DATA_OUT <= DATA_IN(2 DOWNTO 0) & DATA_IN(3);
			WHEN "101"  => DATA_OUT <= DATA_IN(3) & DATA_IN(3 DOWNTO 1);
			WHEN "110"  => DATA_OUT <= DATA_IN(1 DOWNTO 0) & DATA_IN(3 DOWNTO 2);
			WHEN OTHERS => DATA_OUT <= DATA_IN;
		END CASE;
	END PROCESS;
END Hw3Architecture;
